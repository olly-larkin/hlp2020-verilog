module multi_file (
    out
);

output[2:0] out;

CustomCount3 count(out);

endmodule