module multi_file (
    out1
);

output[2:0] out1;

CustomCount3 count(out1);

endmodule